/* -----------------------------------------------
 * Project Name   : DRAC
 * File           : branch_predictor.sv
 * Organization   : Barcelona Supercomputing Center
 * Author(s)      : Victor Soria
 * Email(s)       : victor.soria@bsc.es
 * References     : 
 * -----------------------------------------------
 * Revision History
 *  Revision   | Author    | Commit | Description
 *  0.1        | Victor.SP | 
 * -----------------------------------------------
 */
 
//`default_nettype none
import drac_pkg::*;
import riscv_pkg::*;
 
 // Number of entries of the is branch predictor.
localparam NUM_IS_BRANCH_ENTRIES = 1024; 

// Tags stored in is_branch_table
typedef logic [27:0] tag;
typedef reg   [27:0] tag_reg;

 
/* Top view of the branch predictor module
 * 
 * Describes the different components of the branch prediction unit and 
 * how they are connected. It is composed by Bimodal Predictor and Return
 * Addres Stack.
 */
module branch_predictor(
    input wire           rstn_i,                        // Negative reset input signal
    input wire           clk_i,                         // Clock input signal
    input addrPC_t       pc_fetch_i,                    // Program counter value at Fetch Stage
    input addrPC_t       pc_execution_i,                // Program counter at Execution Stage
    input addrPC_t        branch_addr_result_exec_i,     // Address generated by branch in Execution Stage (for RAS push as well)
    input wire           branch_taken_result_exec_i,    // Taken or not taken branch result in Execution Stage
    input wire           is_branch_EX_i,                // The instruction in the Execution Stage is a branch
    input wire           push_return_address_i,         // Push return_addrPC_to_store_i in RAS 
    input wire           pop_return_address_i,          // Pop the first addr of the RAS to read

    output logic         branch_predict_is_branch_o,    // Bit that encodes if the instruction being fetched is a branch
    output logic         branch_predict_taken_o,        // Bit that encodes branch taken '1' or not '0'
    output addrPC_t      branch_predict_addr_o          // Address predicted to jump
);

////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////
/////////// Declaration of local signals and modules                                               /////////////////////
////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////
                
wire            bimodal_predict_taken;
addrPC_t        bimodal_predict_addr;
tag_reg         is_branch_tag;
addrPC_t        ras_addr;
wire            use_bimodal;
wire            is_branch_prediction;
                
// Instatiation of bimodal predictor
bimodal_predictor bimodal_predictor_inst(
    .rstn_i (rstn_i),
    .clk_i (clk_i),
    .pc_fetch_i (pc_fetch_i),
    .pc_execution_i (pc_execution_i),
    .branch_addr_result_exec_i (branch_addr_result_exec_i),
    .branch_taken_result_exec_i (branch_taken_result_exec_i),
    .is_branch_EX_i (is_branch_EX_i),
    .bimodal_predict_taken_o (bimodal_predict_taken),
    .bimodal_predict_addr_o (bimodal_predict_addr)
);

////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////
/////////// Instantiation of is branch predictor                                                   /////////////////////
////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////

`ifndef SRAM_MEMORIES
    logic [27 : 0] is_branch_table [0 : NUM_IS_BRANCH_ENTRIES-1]; 

    always_ff @(negedge clk_i, negedge rstn_i) 
    begin
        if(~rstn_i) begin
            is_branch_tag <= 'h0;
        end else begin
            is_branch_tag <= is_branch_table[pc_fetch_i[11:2]];
        end
    end
    
    always_ff @(posedge clk_i) 
    begin
         if(is_branch_EX_i) begin
            is_branch_table[pc_execution_i[11:2]] <= pc_execution_i[39:12];
        end
    end


`else  // If SRAM memories are used

    TSDN65LPA1024X28M4S BIPCArray (
        .AA  (write_address) ,
        .DA  (aux_write_data) ,
        .BWEBA  (28'b0) ,
        .WEBA  (!write) ,
        .CEBA  (1'b0) ,
        .CLKA  (clk) ,
        .AB  (aux_read_address) ,
        .DB  (28'b0) ,
        .BWEBB  ({28{1'b1}}) ,
        .WEBB  (1'b1) ,
        .CEBB  (Stall) ,
        .CLKB  (clk) ,
        .QB  (aux_read_data)
    ); // QA output left unconnected

`endif

/*
// Instatiation of RAS.
return_address_stack return_address_stack_inst(
    .rstn_i(rstn_i),
    .clk_i (clk_i),
    .pc_execution_i (pc_execution_i),
    .push_i(push_return_address_i),
    .pop_i(pop_return_address_i),
    .return_address_o(ras_addr)
);*/

assign use_bimodal = 1'b1; // !pop
assign is_branch_prediction = (is_branch_tag == pc_fetch_i[39:12]);


// MUX that decides wheter the predicted address comes from Bimodal or RAS
assign branch_predict_addr_o = (use_bimodal) ? bimodal_predict_addr : ras_addr;

// MUX that decides wheter the branch prediction is comes from Bimodal or RAS
assign branch_predict_taken_o = (use_bimodal) ? bimodal_predict_taken : 1'b1;

// MUX that decides whteter the fetched instruction is a branch or not
assign branch_predict_is_branch_o = (use_bimodal) ? is_branch_prediction : 1'b0;

endmodule
