/* -----------------------------------------------
 * Project Name   : DRAC
 * File           : bimodal_predictor.sv
 * Organization   : Barcelona Supercomputing Center
 * Author(s)      : Victor Soria
 * Email(s)       : victor.soria@bsc.es
 * References     : 
 * -----------------------------------------------
 * Revision History
 *  Revision   | Author    | Commit | Description
 *  0.1        | Victor.SP | 
 * -----------------------------------------------
 */

import drac_pkg::*;
import riscv_pkg::*;

// Length of the bimodal index register
localparam _LENGTH_BIMODAL_INDEX_  = 10;

// Number of entries of the bimodal predictor, must be 2^(_LENGTH_BIMODAL_INDEX_)
localparam _NUM_BIMODAL_ENTRIES_ = 1024;

// Number of bits used for encoding the state of predictor state machine
localparam _BITS_BIMODAL_STATE_MACHINE_ = 2;

// Initial state of the predictor state machine
localparam _INITIAL_STATE_BIMODAL_ = 2'b10;

 
 /* Bimodal branch predictor implementation
  *
  *
  */
module bimodal_predictor(
    input               clk_i,                         // Clock input signal
    input   addrPC_t    pc_fetch_i,                    // Program counter value at Fetch Stage
    input   addrPC_t    pc_execution_i,                // Program counter at Execution Stage
    input   addrPC_t    branch_addr_result_exec_i,     // Address generated by branch in Execution Stage
    input               branch_taken_result_exec_i,    // Taken or not taken branch in Execution Stage
    input               is_branch_EX_i,                // The instruction in the Execution Stage is a branch
    output              bimodal_predict_taken_o,       // Bit that encodes branch taken '1' or not '0'
    output  addrPC_t    bimodal_predict_addr_o         // Address predicted to jump
);

reg [_BITS_BIMODAL_STATE_MACHINE_-1:0] new_state_to_pht;
reg [_BITS_BIMODAL_STATE_MACHINE_-1:0] readed_state_pht;
reg [1:0] past_state_pht;

`ifndef SRAM_MEMORIES

    // Creates an array of _NUM_BIMODAL_ENTRIES_ registers of _BITS_BIMODAL_STATE_MACHINE_ length
    // This array stores 1024 states machines for predicting the branches

    reg [_BITS_BIMODAL_STATE_MACHINE_ -1:0] pattern_history_table [0:_NUM_BIMODAL_ENTRIES_ -1]; 
    reg [63:0] branch_target_buffer [0:_NUM_BIMODAL_ENTRIES_-1];

    
    `ifndef SYNTHESIS
        // Initialize all the entries of the pattern history table with the initial state
        integer i;
        initial 
        begin for(i = 0; i < _NUM_BIMODAL_ENTRIES_ ; i = i + 1) begin
                pattern_history_table[i] = _INITIAL_STATE_BIMODAL_;
                branch_target_buffer[i] = 64'h0;
              end
        end
    `endif


    // Read pattern history table at addres pc_fetch_i
    always@(negedge clk_i)
    begin
        readed_state_pht <= pattern_history_table[pc_fetch_i[MOST_SIGNIFICATIVE_INDEX_BIT_BP:LEAST_SIGNIFICATIVE_INDEX_BIT_BP]];
        past_state_pht <= pattern_history_table[pc_execution_i[MOST_SIGNIFICATIVE_INDEX_BIT_BP:LEAST_SIGNIFICATIVE_INDEX_BIT_BP]];
        bimodal_predict_addr_o <= branch_target_buffer[pc_fetch_i[MOST_SIGNIFICATIVE_INDEX_BIT_BP:LEAST_SIGNIFICATIVE_INDEX_BIT_BP]];
    end
   
    always_comb begin
        if (past_state_pht == 2'b00 && branch_taken_result_exec_i == 1'b0)
            new_state_to_pht = 2'b00;
        else if (past_state_pht == 2'b11 && branch_taken_result_exec_i == 1'b1)
            new_state_to_pht = 2'b11;
        else if (branch_taken_result_exec_i == 1'b1)
            new_state_to_pht = past_state_pht + 2'b01;
        else
            new_state_to_pht = past_state_pht - 2'b01;
    end


    // Write pattern history table at addres pc_fetch_i
    always@(posedge clk_i)
    begin 
        if(is_branch_EX_i) 
            pattern_history_table[pc_execution_i[MOST_SIGNIFICATIVE_INDEX_BIT_BP:LEAST_SIGNIFICATIVE_INDEX_BIT_BP]] <= new_state_to_pht;
            branch_target_buffer[pc_execution_i[MOST_SIGNIFICATIVE_INDEX_BIT_BP:LEAST_SIGNIFICATIVE_INDEX_BIT_BP]] <= branch_addr_result_exec_i;
    end 
    
    // If state is 00 or 01 predict not taken, if 10 or 11 predict taken
    assign bimodal_predict_taken_o = readed_state_pht[1];
 


    
`else // If SRAM memories are used

    // Creates a SRAM table with 1024 entries of 2 bits. It is NOT parametrical.
    // The table has 2 read/write ports
    // This table stores the states machines for predicting the branches

    // Port A: Write; Port B: Read
    TSDN65LPA1024X2M4S pattern_history_table (
        .AA  (pc_execution_i[MOST_SIGNIFICATIVE_INDEX_BIT_BP:LEAST_SIGNIFICATIVE_INDEX_BIT_BP]) ,     // Address port A
        .DA  (new_state_to_pht) ,    // Data write port A
        .BWEBA  (2'b0) ,             //
        .WEBA  (!write) ,            //
        .CEBA  (1'b0) ,              // 
        .CLKA  (clk_i) ,               // Clock port B
        .AB  (aux_read_address) ,    // Address port B
        .DB  (2'b0) ,                // Data port B
        .BWEBB  (2'b11) ,            //
        .WEBB  (1'b1) ,              //
        .CEBB  (Stall) ,             //
        .CLKB  (clk_i) ,             // Clock port B
        .QB  (aux_read_data)         // Read port B
    ); // QA output left unconnected

`endif

endmodule
