//Write a nice header
