`ifndef TEST_CONSTS_H
  `define TEST_CONSTS_H

	`define N_TESTS            'd100  // Number of random reads in test
	`define ADDR_MIN           'd0   // minimum addr range for read operations
	`define ADDR_MAX           'd524287 // maximum addr range for read operations

`endif
