/*
 * Copyright 2025 BSC*
 * *Barcelona Supercomputing Center (BSC)
 * 
 * SPDX-License-Identifier: Apache-2.0 WITH SHL-2.1
 * 
 * Licensed under the Solderpad Hardware License v 2.1 (the “License”); you
 * may not use this file except in compliance with the License, or, at your
 * option, the Apache License version 2.0. You may obtain a copy of the
 * License at
 * 
 * https://solderpad.org/licenses/SHL-2.1/
 * 
 * Unless required by applicable law or agreed to in writing, any work
 * distributed under the License is distributed on an “AS IS” BASIS, WITHOUT
 * WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied. See the
 * License for the specific language governing permissions and limitations
 * under the License.
 */
 
 /* Bimodal branch predictor implementation
  *
  *
  */
module bimodal_predictor
    import drac_pkg::*;
    import riscv_pkg::*;
(
    input   logic       clk_i,                         // Clock input signal
    input   logic       rstn_i,                        // reset input signal
    input   addrPC_t    pc_fetch_i,                    // Program counter value at Fetch Stage
    input   addrPC_t    pc_execution_i,                // Program counter at Execution Stage
    input   addrPC_t    branch_addr_result_exec_i,     // Address generated by branch in Execution Stage
    input   logic       branch_taken_result_exec_i,    // Taken or not taken branch in Execution Stage
    input   logic       is_branch_EX_i,                // The instruction in the Execution Stage is a branch
    output  logic       bimodal_predict_taken_o,       // Bit that encodes branch taken '1' or not '0'
    output  addrPC_t    bimodal_predict_addr_o         // Address predicted to jump
);

// Length of the bimodal index register
localparam _LENGTH_BIMODAL_INDEX_  = 7;
// Number of entries of the bimodal predictor, must be 2^(_LENGTH_BIMODAL_INDEX_)
localparam _NUM_BIMODAL_ENTRIES_ = 2**_LENGTH_BIMODAL_INDEX_;
// Number of bits used for encoding the state of predictor state machine
localparam _BITS_BIMODAL_STATE_MACHINE_ = 2;

function [_BITS_BIMODAL_STATE_MACHINE_-1:0] trunc_bp_sum(input [_BITS_BIMODAL_STATE_MACHINE_:0] val_in);
    trunc_bp_sum = val_in[_BITS_BIMODAL_STATE_MACHINE_-1:0];
endfunction

logic [_BITS_BIMODAL_STATE_MACHINE_-1:0] new_state_to_pht;
logic [_BITS_BIMODAL_STATE_MACHINE_-1:0] readed_state_pht;
logic [1:0] past_state_pht;

    // Creates an array of _NUM_BIMODAL_ENTRIES_ registers of _BITS_BIMODAL_STATE_MACHINE_ length
    // This array stores 1024 states machines for predicting the branches

    reg [_BITS_BIMODAL_STATE_MACHINE_ -1:0] pattern_history_table [_NUM_BIMODAL_ENTRIES_-1:0]; 
    // We need to store the PHY_VIRT_MAX_ADDR_SIZE + 1 bits in order to perform properly the sign extension 
    reg [PHY_VIRT_MAX_ADDR_SIZE:0] branch_target_buffer [_NUM_BIMODAL_ENTRIES_-1:0];

    // Read pattern history table at addres pc_fetch_i
    logic [PHY_VIRT_MAX_ADDR_SIZE:0] short_pred_addr;
    always_comb
    begin
        readed_state_pht = pattern_history_table[pc_fetch_i[MOST_SIGNIFICATIVE_INDEX_BIT_BP:LEAST_SIGNIFICATIVE_INDEX_BIT_BP]];
        past_state_pht = pattern_history_table[pc_execution_i[MOST_SIGNIFICATIVE_INDEX_BIT_BP:LEAST_SIGNIFICATIVE_INDEX_BIT_BP]];
        short_pred_addr = branch_target_buffer[pc_fetch_i[MOST_SIGNIFICATIVE_INDEX_BIT_BP:LEAST_SIGNIFICATIVE_INDEX_BIT_BP]];
        bimodal_predict_addr_o = { {(XLEN-PHY_VIRT_MAX_ADDR_SIZE-1){short_pred_addr[PHY_VIRT_MAX_ADDR_SIZE]}}, short_pred_addr};
    end
   
    always_comb begin
        if ((past_state_pht == 2'b00) && (branch_taken_result_exec_i == 1'b0))
            new_state_to_pht = 2'b00;
        else if ((past_state_pht == 2'b11) && (branch_taken_result_exec_i == 1'b1))
            new_state_to_pht = 2'b11;
        else if (branch_taken_result_exec_i == 1'b1)
            new_state_to_pht = trunc_bp_sum(past_state_pht + 2'b01);
        else
            new_state_to_pht = trunc_bp_sum(past_state_pht - 2'b01);
    end


    // Write pattern history table at addres pc_fetch_i
    always_ff @(posedge clk_i or negedge rstn_i ) begin 
		if (~rstn_i) begin
			for(integer i = 0; i < _NUM_BIMODAL_ENTRIES_ ; i = i + 1) begin
				pattern_history_table[i] <= 2'b01;
                branch_target_buffer[i] <= 'h0;
			end
        end else if(is_branch_EX_i) begin 
            pattern_history_table[pc_execution_i[MOST_SIGNIFICATIVE_INDEX_BIT_BP:LEAST_SIGNIFICATIVE_INDEX_BIT_BP]] <= new_state_to_pht;
            branch_target_buffer[pc_execution_i[MOST_SIGNIFICATIVE_INDEX_BIT_BP:LEAST_SIGNIFICATIVE_INDEX_BIT_BP]] <= branch_addr_result_exec_i[PHY_VIRT_MAX_ADDR_SIZE:0];
		end
    end    
    // If state is 00 or 01 predict not taken, if 10 or 11 predict taken
    assign bimodal_predict_taken_o = readed_state_pht[1];

endmodule
