`ifndef TEST_CONSTS_H
  `define TEST_CONSTS_H

  parameter N_TESTS  = 'd100;  // Number of random reads in test
  parameter ADDR_MIN = 'd0;   // minimum addr range for read operations
  parameter ADDR_MAX = 'd524287; // maximum addr range for read operations
  

`endif
