//DRAC
